module ALU_DUT();
//input
 reg  signed [15:0] A, B;
 reg signed [2:0] OP;
 //output
 wire  signed [31:0] ALU_OUTPUT;
 //simulation
 initial
 begin
      //        Addition
 // 16'b111100 + 16'b1111 = 32'1001011 (75)
  OP = 3'b000 ; A = 60 ; B = 15 ; #10;
 // 0 + 4000 = 4000
  OP = 3'b000 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 + 8000 = 16000
  OP = 3'b000 ; A = 16'd8000 ; B = 16'd8000 ; #10;
//3000 + 9000 = 12000
  OP = 3'b000 ; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 + 40 = -40
  OP = 3'b000 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 + (-21) =-63
  OP = 3'b000 ; A = -16'd42 ; B = -16'd21 ; #10;


         //        subtraction
// 16'b111100 - 16'b1111 = 32'101101 (45)
  OP = 3'b001 ; A = 60 ; B = 15 ; #10;
// 0 - 4000 = -4000
  OP = 3'b001 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 - 8000 = 0
  OP = 3'b001 ; A = 16'd8000 ; B = 16'd8000 ; #10;
// 3000 - 9000 = -6000
  OP = 3'b001 ; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 - 40 = -120
  OP = 3'b001 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 - (-21) =-21
  OP = 3'b001 ; A = -16'd42 ; B = -16'd21 ; #10;


         //        Multiplication
// 16'b111100 * 16'b1111 = 32'1110000100 (900)
  OP = 3'b010 ; A = 60 ; B = 15 ; #10;
//0 * 4000 = 0
  OP = 3'b010 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 * 8000 = 64000000
  OP = 3'b010 ; A = 16'd8000 ; B = 16'd8000 ; #10;
// 3000 * 9000 = 27000000
  OP = 3'b010 ; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 * 40 = -3200
  OP = 3'b010 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 * (-21) = 882
  OP = 3'b010 ; A = -16'd42 ; B = -16'd21 ; #10;


         //        Division
// 16'b111100 / 16'b1111 = 32'b100 (4)
  OP = 3'b011 ; A = 60 ; B = 15 ; #10;
//0 / 4000 = 0
  OP = 3'b011 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 / 8000 = 1 
  OP = 3'b011 ; A = 16'd8000 ; B = 16'd8000 ; #10;
// 3000 / 9000 = 0 (INTEGER)
  OP = 3'b011; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 / 40 = -2
  OP = 3'b011 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 / (-21) =2
  OP = 3'b011 ; A = -16'd42 ; B = -16'd21 ; #10;




        //        OR Gate
// 16'b111100 | 16'b1111 = 32'1111111
  OP = 3'b100 ; A = 60 ; B = 15 ; #10;
// 0 OR 4000 
  OP = 3'b100 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 OR 8000 
  OP = 3'b100 ; A = 16'd8000 ; B = 16'd8000 ; #10;
// 3000 OR 9000 
  OP = 3'b100 ; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 OR 40 
  OP = 3'b100 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 OR (-21)  
  OP = 3'b100 ; A = -16'd42 ; B = -16'd21 ; #10;


         //        AND Gate
// 16'b111100 & 16'b1111 = 32'1100
  OP = 3'b101 ; A = 60 ; B = 15 ; #10;
// 0 and 4000
  OP = 3'b101 ; A = 16'd0 ; B = 16'd4000 ; #10;
// 8000 AND 8000
  OP = 3'b101 ; A = 16'd8000 ; B = 16'd8000 ; #10;
// 3000 AND 9000 
  OP = 3'b101 ; A = 16'd3000 ; B = 16'd9000 ; #10;
//-80 AND 40
  OP = 3'b101 ; A = -16'd80 ; B = 16'd40 ; #10;
//-42 AND (-21) 
  OP = 3'b101 ; A = -16'd42 ; B = -16'd21 ; #10;


        //        not A
// not A 
  OP = 3'b110 ; A = 60 ; B = 15 ; #10;
  OP = 3'b110 ; A = 16'd0 ; B = 16'd4000 ; #10;
  OP = 3'b110 ; A = 16'd8000 ; B = 16'd8000 ; #10;
  OP = 3'b110 ; A = 16'd3000 ; B = 16'd9000 ; #10;
  OP = 3'b110 ; A = -16'd80 ; B = 16'd40 ; #10;
  OP = 3'b110 ; A = -16'd42 ; B = -16'd21 ; #10;

         //        not B
  OP = 3'b111 ; A = 60 ; B = 15 ; #10;
  OP = 3'b111 ; A = 16'd0 ; B = 16'd4000 ; #10;
  OP = 3'b111 ; A = 16'd8000 ; B = 16'd8000 ; #10;
  OP = 3'b111 ; A = 16'd3000 ; B = 16'd9000 ; #10;
  OP = 3'b111 ; A = -16'd80 ; B = 16'd40 ; #10;
  OP = 3'b111 ; A = -16'd42 ; B = -16'd21 ; #10;
 end
 ALU ALU1(A, B, OP, ALU_OUTPUT);
initial begin
$display("    B      A           output   ");
$monitor(" %b    %b = %b ",A,   B,   ALU_OUTPUT);
end 
endmodule 
